*Simple n-input OTA


.param Wtail_currrent = 
.param Ltail_current = 

.param WM6 = 
.param LM6 = 

.param W5 =
.param L5 =

.param W4 =
.param L4 =

.param W3 = 
.param L3 = 

.subckt simple_nmos ninp ninn noutp noutn nbias1 nbias2 ndd nss

X_M6a out_p b5 vdd vdd pmos w=WM6 L=LM6
X_M6b out_n b5 vdd vdd pmos w=WM6 L=LM6

X_M5a pout b4 out_p vdd pmos w=W5 L=L5
X_M5b nout b4 out_n vdd pmos w=W5 L=L5

X_M4a pout b3 m4a_source nss nmos w=W4 L=L4
X_M4b nout b3 m4b_source nss nmos w=W4 L=L4

X_M3a m4a_source b2 nss nss pmos w=W3 L=L3
X_M3b m4b_source b2 nss nss pmos w=W3 L=L3

X_inpPair_p out_p inp_n tail_node nss nmos w=Winp_pair l=Linp_pair
X_inpPair_n out_n inp_p tail_node nss nmos w=Winp_pair l=Linp_pair


X_tailCurrentSource tail_node nbias1 nss nss nmos w=Wtail_current l=Ltail_current

.ends simple_nmos
